module nor_gate(
input a,b,
output y);
nor n1(y,a,b);
endmodule

