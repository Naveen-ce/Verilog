module and_gate
