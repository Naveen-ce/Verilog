module not_gate(
input a,
output y);
not n1(y,a);
endmodule
