module xnor_gate(
input a,b,
output y);
xnor x1(y,a,b);
endmodule
