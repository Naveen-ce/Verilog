module or_gate(
input a,b,
output y);
or o1(y,a,b);
endmodule
