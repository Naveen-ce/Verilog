module divide;
integer b;
initial
begin
b=-‘d 12/3;
$display("b=%d",b);
end
endmodule
