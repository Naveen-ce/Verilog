module async_up_counter(
input
